module aig_mix_5_vl5(
    input [127:0] in,
    output [63:0] out
);

// Mixed AIG logic with various patterns
wire [255:0] internal;

assign internal[0] = in[0] & in[0];
assign internal[1] = in[7] | in[11];
assign internal[2] = in[14] ^ in[22];
assign internal[3] = ~(in[21] & in[33] & in[39]);
assign internal[4] = in[28] & in[44];
assign internal[5] = in[35] | in[55];
assign internal[6] = in[42] ^ in[66];
assign internal[7] = ~(in[49] & in[77] & in[91]);
assign internal[8] = in[56] & in[88];
assign internal[9] = in[63] | in[99];
assign internal[10] = in[70] ^ in[110];
assign internal[11] = ~(in[77] & in[121] & in[15]);
assign internal[12] = in[84] & in[4];
assign internal[13] = in[91] | in[15];
assign internal[14] = in[98] ^ in[26];
assign internal[15] = ~(in[105] & in[37] & in[67]);
assign internal[16] = in[112] & in[48];
assign internal[17] = in[119] | in[59];
assign internal[18] = in[126] ^ in[70];
assign internal[19] = ~(in[5] & in[81] & in[119]);
assign internal[20] = in[12] & in[92];
assign internal[21] = in[19] | in[103];
assign internal[22] = in[26] ^ in[114];
assign internal[23] = ~(in[33] & in[125] & in[43]);
assign internal[24] = in[40] & in[8];
assign internal[25] = in[47] | in[19];
assign internal[26] = in[54] ^ in[30];
assign internal[27] = ~(in[61] & in[41] & in[95]);
assign internal[28] = in[68] & in[52];
assign internal[29] = in[75] | in[63];
assign internal[30] = in[82] ^ in[74];
assign internal[31] = ~(in[89] & in[85] & in[19]);
assign internal[32] = in[96] & in[96];
assign internal[33] = in[103] | in[107];
assign internal[34] = in[110] ^ in[118];
assign internal[35] = ~(in[117] & in[1] & in[71]);
assign internal[36] = in[124] & in[12];
assign internal[37] = in[3] | in[23];
assign internal[38] = in[10] ^ in[34];
assign internal[39] = ~(in[17] & in[45] & in[123]);
assign internal[40] = in[24] & in[56];
assign internal[41] = in[31] | in[67];
assign internal[42] = in[38] ^ in[78];
assign internal[43] = ~(in[45] & in[89] & in[47]);
assign internal[44] = in[52] & in[100];
assign internal[45] = in[59] | in[111];
assign internal[46] = in[66] ^ in[122];
assign internal[47] = ~(in[73] & in[5] & in[99]);
assign internal[48] = in[80] & in[16];
assign internal[49] = in[87] | in[27];
assign internal[50] = in[94] ^ in[38];
assign internal[51] = ~(in[101] & in[49] & in[23]);
assign internal[52] = in[108] & in[60];
assign internal[53] = in[115] | in[71];
assign internal[54] = in[122] ^ in[82];
assign internal[55] = ~(in[1] & in[93] & in[75]);
assign internal[56] = in[8] & in[104];
assign internal[57] = in[15] | in[115];
assign internal[58] = in[22] ^ in[126];
assign internal[59] = ~(in[29] & in[9] & in[127]);
assign internal[60] = in[36] & in[20];
assign internal[61] = in[43] | in[31];
assign internal[62] = in[50] ^ in[42];
assign internal[63] = ~(in[57] & in[53] & in[51]);
assign internal[64] = in[64] & in[64];
assign internal[65] = in[71] | in[75];
assign internal[66] = in[78] ^ in[86];
assign internal[67] = ~(in[85] & in[97] & in[103]);
assign internal[68] = in[92] & in[108];
assign internal[69] = in[99] | in[119];
assign internal[70] = in[106] ^ in[2];
assign internal[71] = ~(in[113] & in[13] & in[27]);
assign internal[72] = in[120] & in[24];
assign internal[73] = in[127] | in[35];
assign internal[74] = in[6] ^ in[46];
assign internal[75] = ~(in[13] & in[57] & in[79]);
assign internal[76] = in[20] & in[68];
assign internal[77] = in[27] | in[79];
assign internal[78] = in[34] ^ in[90];
assign internal[79] = ~(in[41] & in[101] & in[3]);
assign internal[80] = in[48] & in[112];
assign internal[81] = in[55] | in[123];
assign internal[82] = in[62] ^ in[6];
assign internal[83] = ~(in[69] & in[17] & in[55]);
assign internal[84] = in[76] & in[28];
assign internal[85] = in[83] | in[39];
assign internal[86] = in[90] ^ in[50];
assign internal[87] = ~(in[97] & in[61] & in[107]);
assign internal[88] = in[104] & in[72];
assign internal[89] = in[111] | in[83];
assign internal[90] = in[118] ^ in[94];
assign internal[91] = ~(in[125] & in[105] & in[31]);
assign internal[92] = in[4] & in[116];
assign internal[93] = in[11] | in[127];
assign internal[94] = in[18] ^ in[10];
assign internal[95] = ~(in[25] & in[21] & in[83]);
assign internal[96] = in[32] & in[32];
assign internal[97] = in[39] | in[43];
assign internal[98] = in[46] ^ in[54];
assign internal[99] = ~(in[53] & in[65] & in[7]);
assign internal[100] = in[60] & in[76];
assign internal[101] = in[67] | in[87];
assign internal[102] = in[74] ^ in[98];
assign internal[103] = ~(in[81] & in[109] & in[59]);
assign internal[104] = in[88] & in[120];
assign internal[105] = in[95] | in[3];
assign internal[106] = in[102] ^ in[14];
assign internal[107] = ~(in[109] & in[25] & in[111]);
assign internal[108] = in[116] & in[36];
assign internal[109] = in[123] | in[47];
assign internal[110] = in[2] ^ in[58];
assign internal[111] = ~(in[9] & in[69] & in[35]);
assign internal[112] = in[16] & in[80];
assign internal[113] = in[23] | in[91];
assign internal[114] = in[30] ^ in[102];
assign internal[115] = ~(in[37] & in[113] & in[87]);
assign internal[116] = in[44] & in[124];
assign internal[117] = in[51] | in[7];
assign internal[118] = in[58] ^ in[18];
assign internal[119] = ~(in[65] & in[29] & in[11]);
assign internal[120] = in[72] & in[40];
assign internal[121] = in[79] | in[51];
assign internal[122] = in[86] ^ in[62];
assign internal[123] = ~(in[93] & in[73] & in[63]);
assign internal[124] = in[100] & in[84];
assign internal[125] = in[107] | in[95];
assign internal[126] = in[114] ^ in[106];
assign internal[127] = ~(in[121] & in[117] & in[115]);
assign internal[128] = in[0] & in[0];
assign internal[129] = in[7] | in[11];
assign internal[130] = in[14] ^ in[22];
assign internal[131] = ~(in[21] & in[33] & in[39]);
assign internal[132] = in[28] & in[44];
assign internal[133] = in[35] | in[55];
assign internal[134] = in[42] ^ in[66];
assign internal[135] = ~(in[49] & in[77] & in[91]);
assign internal[136] = in[56] & in[88];
assign internal[137] = in[63] | in[99];
assign internal[138] = in[70] ^ in[110];
assign internal[139] = ~(in[77] & in[121] & in[15]);
assign internal[140] = in[84] & in[4];
assign internal[141] = in[91] | in[15];
assign internal[142] = in[98] ^ in[26];
assign internal[143] = ~(in[105] & in[37] & in[67]);
assign internal[144] = in[112] & in[48];
assign internal[145] = in[119] | in[59];
assign internal[146] = in[126] ^ in[70];
assign internal[147] = ~(in[5] & in[81] & in[119]);
assign internal[148] = in[12] & in[92];
assign internal[149] = in[19] | in[103];
assign internal[150] = in[26] ^ in[114];
assign internal[151] = ~(in[33] & in[125] & in[43]);
assign internal[152] = in[40] & in[8];
assign internal[153] = in[47] | in[19];
assign internal[154] = in[54] ^ in[30];
assign internal[155] = ~(in[61] & in[41] & in[95]);
assign internal[156] = in[68] & in[52];
assign internal[157] = in[75] | in[63];
assign internal[158] = in[82] ^ in[74];
assign internal[159] = ~(in[89] & in[85] & in[19]);
assign internal[160] = in[96] & in[96];
assign internal[161] = in[103] | in[107];
assign internal[162] = in[110] ^ in[118];
assign internal[163] = ~(in[117] & in[1] & in[71]);
assign internal[164] = in[124] & in[12];
assign internal[165] = in[3] | in[23];
assign internal[166] = in[10] ^ in[34];
assign internal[167] = ~(in[17] & in[45] & in[123]);
assign internal[168] = in[24] & in[56];
assign internal[169] = in[31] | in[67];
assign internal[170] = in[38] ^ in[78];
assign internal[171] = ~(in[45] & in[89] & in[47]);
assign internal[172] = in[52] & in[100];
assign internal[173] = in[59] | in[111];
assign internal[174] = in[66] ^ in[122];
assign internal[175] = ~(in[73] & in[5] & in[99]);
assign internal[176] = in[80] & in[16];
assign internal[177] = in[87] | in[27];
assign internal[178] = in[94] ^ in[38];
assign internal[179] = ~(in[101] & in[49] & in[23]);
assign internal[180] = in[108] & in[60];
assign internal[181] = in[115] | in[71];
assign internal[182] = in[122] ^ in[82];
assign internal[183] = ~(in[1] & in[93] & in[75]);
assign internal[184] = in[8] & in[104];
assign internal[185] = in[15] | in[115];
assign internal[186] = in[22] ^ in[126];
assign internal[187] = ~(in[29] & in[9] & in[127]);
assign internal[188] = in[36] & in[20];
assign internal[189] = in[43] | in[31];
assign internal[190] = in[50] ^ in[42];
assign internal[191] = ~(in[57] & in[53] & in[51]);
assign internal[192] = in[64] & in[64];
assign internal[193] = in[71] | in[75];
assign internal[194] = in[78] ^ in[86];
assign internal[195] = ~(in[85] & in[97] & in[103]);
assign internal[196] = in[92] & in[108];
assign internal[197] = in[99] | in[119];
assign internal[198] = in[106] ^ in[2];
assign internal[199] = ~(in[113] & in[13] & in[27]);
assign internal[200] = in[120] & in[24];
assign internal[201] = in[127] | in[35];
assign internal[202] = in[6] ^ in[46];
assign internal[203] = ~(in[13] & in[57] & in[79]);
assign internal[204] = in[20] & in[68];
assign internal[205] = in[27] | in[79];
assign internal[206] = in[34] ^ in[90];
assign internal[207] = ~(in[41] & in[101] & in[3]);
assign internal[208] = in[48] & in[112];
assign internal[209] = in[55] | in[123];
assign internal[210] = in[62] ^ in[6];
assign internal[211] = ~(in[69] & in[17] & in[55]);
assign internal[212] = in[76] & in[28];
assign internal[213] = in[83] | in[39];
assign internal[214] = in[90] ^ in[50];
assign internal[215] = ~(in[97] & in[61] & in[107]);
assign internal[216] = in[104] & in[72];
assign internal[217] = in[111] | in[83];
assign internal[218] = in[118] ^ in[94];
assign internal[219] = ~(in[125] & in[105] & in[31]);
assign internal[220] = in[4] & in[116];
assign internal[221] = in[11] | in[127];
assign internal[222] = in[18] ^ in[10];
assign internal[223] = ~(in[25] & in[21] & in[83]);
assign internal[224] = in[32] & in[32];
assign internal[225] = in[39] | in[43];
assign internal[226] = in[46] ^ in[54];
assign internal[227] = ~(in[53] & in[65] & in[7]);
assign internal[228] = in[60] & in[76];
assign internal[229] = in[67] | in[87];
assign internal[230] = in[74] ^ in[98];
assign internal[231] = ~(in[81] & in[109] & in[59]);
assign internal[232] = in[88] & in[120];
assign internal[233] = in[95] | in[3];
assign internal[234] = in[102] ^ in[14];
assign internal[235] = ~(in[109] & in[25] & in[111]);
assign internal[236] = in[116] & in[36];
assign internal[237] = in[123] | in[47];
assign internal[238] = in[2] ^ in[58];
assign internal[239] = ~(in[9] & in[69] & in[35]);
assign internal[240] = in[16] & in[80];
assign internal[241] = in[23] | in[91];
assign internal[242] = in[30] ^ in[102];
assign internal[243] = ~(in[37] & in[113] & in[87]);
assign internal[244] = in[44] & in[124];
assign internal[245] = in[51] | in[7];
assign internal[246] = in[58] ^ in[18];
assign internal[247] = ~(in[65] & in[29] & in[11]);
assign internal[248] = in[72] & in[40];
assign internal[249] = in[79] | in[51];
assign internal[250] = in[86] ^ in[62];
assign internal[251] = ~(in[93] & in[73] & in[63]);
assign internal[252] = in[100] & in[84];
assign internal[253] = in[107] | in[95];
assign internal[254] = in[114] ^ in[106];
assign internal[255] = ~(in[121] & in[117] & in[115]);

assign out[0] = internal[0] & internal[0];
assign out[1] = internal[3] | internal[5];
assign out[2] = internal[6] ^ internal[10] ^ internal[14];
assign out[3] = internal[9] & internal[15];
assign out[4] = internal[12] | internal[20];
assign out[5] = internal[15] ^ internal[25] ^ internal[35];
assign out[6] = internal[18] & internal[30];
assign out[7] = internal[21] | internal[35];
assign out[8] = internal[24] ^ internal[40] ^ internal[56];
assign out[9] = internal[27] & internal[45];
assign out[10] = internal[30] | internal[50];
assign out[11] = internal[33] ^ internal[55] ^ internal[77];
assign out[12] = internal[36] & internal[60];
assign out[13] = internal[39] | internal[65];
assign out[14] = internal[42] ^ internal[70] ^ internal[98];
assign out[15] = internal[45] & internal[75];
assign out[16] = internal[48] | internal[80];
assign out[17] = internal[51] ^ internal[85] ^ internal[119];
assign out[18] = internal[54] & internal[90];
assign out[19] = internal[57] | internal[95];
assign out[20] = internal[60] ^ internal[100] ^ internal[140];
assign out[21] = internal[63] & internal[105];
assign out[22] = internal[66] | internal[110];
assign out[23] = internal[69] ^ internal[115] ^ internal[161];
assign out[24] = internal[72] & internal[120];
assign out[25] = internal[75] | internal[125];
assign out[26] = internal[78] ^ internal[130] ^ internal[182];
assign out[27] = internal[81] & internal[135];
assign out[28] = internal[84] | internal[140];
assign out[29] = internal[87] ^ internal[145] ^ internal[203];
assign out[30] = internal[90] & internal[150];
assign out[31] = internal[93] | internal[155];
assign out[32] = internal[96] ^ internal[160] ^ internal[224];
assign out[33] = internal[99] & internal[165];
assign out[34] = internal[102] | internal[170];
assign out[35] = internal[105] ^ internal[175] ^ internal[245];
assign out[36] = internal[108] & internal[180];
assign out[37] = internal[111] | internal[185];
assign out[38] = internal[114] ^ internal[190] ^ internal[10];
assign out[39] = internal[117] & internal[195];
assign out[40] = internal[120] | internal[200];
assign out[41] = internal[123] ^ internal[205] ^ internal[31];
assign out[42] = internal[126] & internal[210];
assign out[43] = internal[129] | internal[215];
assign out[44] = internal[132] ^ internal[220] ^ internal[52];
assign out[45] = internal[135] & internal[225];
assign out[46] = internal[138] | internal[230];
assign out[47] = internal[141] ^ internal[235] ^ internal[73];
assign out[48] = internal[144] & internal[240];
assign out[49] = internal[147] | internal[245];
assign out[50] = internal[150] ^ internal[250] ^ internal[94];
assign out[51] = internal[153] & internal[255];
assign out[52] = internal[156] | internal[4];
assign out[53] = internal[159] ^ internal[9] ^ internal[115];
assign out[54] = internal[162] & internal[14];
assign out[55] = internal[165] | internal[19];
assign out[56] = internal[168] ^ internal[24] ^ internal[136];
assign out[57] = internal[171] & internal[29];
assign out[58] = internal[174] | internal[34];
assign out[59] = internal[177] ^ internal[39] ^ internal[157];
assign out[60] = internal[180] & internal[44];
assign out[61] = internal[183] | internal[49];
assign out[62] = internal[186] ^ internal[54] ^ internal[178];
assign out[63] = internal[189] & internal[59];

endmodule