module aig_mix_6_vl6(
    input [143:0] in,
    output [71:0] out
);

// Mixed AIG logic with various patterns
wire [287:0] internal;

assign internal[0] = in[0] & in[0];
assign internal[1] = in[7] | in[11];
assign internal[2] = in[14] ^ in[22];
assign internal[3] = ~(in[21] & in[33] & in[39]);
assign internal[4] = in[28] & in[44];
assign internal[5] = in[35] | in[55];
assign internal[6] = in[42] ^ in[66];
assign internal[7] = ~(in[49] & in[77] & in[91]);
assign internal[8] = in[56] & in[88];
assign internal[9] = in[63] | in[99];
assign internal[10] = in[70] ^ in[110];
assign internal[11] = ~(in[77] & in[121] & in[143]);
assign internal[12] = in[84] & in[132];
assign internal[13] = in[91] | in[143];
assign internal[14] = in[98] ^ in[10];
assign internal[15] = ~(in[105] & in[21] & in[51]);
assign internal[16] = in[112] & in[32];
assign internal[17] = in[119] | in[43];
assign internal[18] = in[126] ^ in[54];
assign internal[19] = ~(in[133] & in[65] & in[103]);
assign internal[20] = in[140] & in[76];
assign internal[21] = in[3] | in[87];
assign internal[22] = in[10] ^ in[98];
assign internal[23] = ~(in[17] & in[109] & in[11]);
assign internal[24] = in[24] & in[120];
assign internal[25] = in[31] | in[131];
assign internal[26] = in[38] ^ in[142];
assign internal[27] = ~(in[45] & in[9] & in[63]);
assign internal[28] = in[52] & in[20];
assign internal[29] = in[59] | in[31];
assign internal[30] = in[66] ^ in[42];
assign internal[31] = ~(in[73] & in[53] & in[115]);
assign internal[32] = in[80] & in[64];
assign internal[33] = in[87] | in[75];
assign internal[34] = in[94] ^ in[86];
assign internal[35] = ~(in[101] & in[97] & in[23]);
assign internal[36] = in[108] & in[108];
assign internal[37] = in[115] | in[119];
assign internal[38] = in[122] ^ in[130];
assign internal[39] = ~(in[129] & in[141] & in[75]);
assign internal[40] = in[136] & in[8];
assign internal[41] = in[143] | in[19];
assign internal[42] = in[6] ^ in[30];
assign internal[43] = ~(in[13] & in[41] & in[127]);
assign internal[44] = in[20] & in[52];
assign internal[45] = in[27] | in[63];
assign internal[46] = in[34] ^ in[74];
assign internal[47] = ~(in[41] & in[85] & in[35]);
assign internal[48] = in[48] & in[96];
assign internal[49] = in[55] | in[107];
assign internal[50] = in[62] ^ in[118];
assign internal[51] = ~(in[69] & in[129] & in[87]);
assign internal[52] = in[76] & in[140];
assign internal[53] = in[83] | in[7];
assign internal[54] = in[90] ^ in[18];
assign internal[55] = ~(in[97] & in[29] & in[139]);
assign internal[56] = in[104] & in[40];
assign internal[57] = in[111] | in[51];
assign internal[58] = in[118] ^ in[62];
assign internal[59] = ~(in[125] & in[73] & in[47]);
assign internal[60] = in[132] & in[84];
assign internal[61] = in[139] | in[95];
assign internal[62] = in[2] ^ in[106];
assign internal[63] = ~(in[9] & in[117] & in[99]);
assign internal[64] = in[16] & in[128];
assign internal[65] = in[23] | in[139];
assign internal[66] = in[30] ^ in[6];
assign internal[67] = ~(in[37] & in[17] & in[7]);
assign internal[68] = in[44] & in[28];
assign internal[69] = in[51] | in[39];
assign internal[70] = in[58] ^ in[50];
assign internal[71] = ~(in[65] & in[61] & in[59]);
assign internal[72] = in[72] & in[72];
assign internal[73] = in[79] | in[83];
assign internal[74] = in[86] ^ in[94];
assign internal[75] = ~(in[93] & in[105] & in[111]);
assign internal[76] = in[100] & in[116];
assign internal[77] = in[107] | in[127];
assign internal[78] = in[114] ^ in[138];
assign internal[79] = ~(in[121] & in[5] & in[19]);
assign internal[80] = in[128] & in[16];
assign internal[81] = in[135] | in[27];
assign internal[82] = in[142] ^ in[38];
assign internal[83] = ~(in[5] & in[49] & in[71]);
assign internal[84] = in[12] & in[60];
assign internal[85] = in[19] | in[71];
assign internal[86] = in[26] ^ in[82];
assign internal[87] = ~(in[33] & in[93] & in[123]);
assign internal[88] = in[40] & in[104];
assign internal[89] = in[47] | in[115];
assign internal[90] = in[54] ^ in[126];
assign internal[91] = ~(in[61] & in[137] & in[31]);
assign internal[92] = in[68] & in[4];
assign internal[93] = in[75] | in[15];
assign internal[94] = in[82] ^ in[26];
assign internal[95] = ~(in[89] & in[37] & in[83]);
assign internal[96] = in[96] & in[48];
assign internal[97] = in[103] | in[59];
assign internal[98] = in[110] ^ in[70];
assign internal[99] = ~(in[117] & in[81] & in[135]);
assign internal[100] = in[124] & in[92];
assign internal[101] = in[131] | in[103];
assign internal[102] = in[138] ^ in[114];
assign internal[103] = ~(in[1] & in[125] & in[43]);
assign internal[104] = in[8] & in[136];
assign internal[105] = in[15] | in[3];
assign internal[106] = in[22] ^ in[14];
assign internal[107] = ~(in[29] & in[25] & in[95]);
assign internal[108] = in[36] & in[36];
assign internal[109] = in[43] | in[47];
assign internal[110] = in[50] ^ in[58];
assign internal[111] = ~(in[57] & in[69] & in[3]);
assign internal[112] = in[64] & in[80];
assign internal[113] = in[71] | in[91];
assign internal[114] = in[78] ^ in[102];
assign internal[115] = ~(in[85] & in[113] & in[55]);
assign internal[116] = in[92] & in[124];
assign internal[117] = in[99] | in[135];
assign internal[118] = in[106] ^ in[2];
assign internal[119] = ~(in[113] & in[13] & in[107]);
assign internal[120] = in[120] & in[24];
assign internal[121] = in[127] | in[35];
assign internal[122] = in[134] ^ in[46];
assign internal[123] = ~(in[141] & in[57] & in[15]);
assign internal[124] = in[4] & in[68];
assign internal[125] = in[11] | in[79];
assign internal[126] = in[18] ^ in[90];
assign internal[127] = ~(in[25] & in[101] & in[67]);
assign internal[128] = in[32] & in[112];
assign internal[129] = in[39] | in[123];
assign internal[130] = in[46] ^ in[134];
assign internal[131] = ~(in[53] & in[1] & in[119]);
assign internal[132] = in[60] & in[12];
assign internal[133] = in[67] | in[23];
assign internal[134] = in[74] ^ in[34];
assign internal[135] = ~(in[81] & in[45] & in[27]);
assign internal[136] = in[88] & in[56];
assign internal[137] = in[95] | in[67];
assign internal[138] = in[102] ^ in[78];
assign internal[139] = ~(in[109] & in[89] & in[79]);
assign internal[140] = in[116] & in[100];
assign internal[141] = in[123] | in[111];
assign internal[142] = in[130] ^ in[122];
assign internal[143] = ~(in[137] & in[133] & in[131]);
assign internal[144] = in[0] & in[0];
assign internal[145] = in[7] | in[11];
assign internal[146] = in[14] ^ in[22];
assign internal[147] = ~(in[21] & in[33] & in[39]);
assign internal[148] = in[28] & in[44];
assign internal[149] = in[35] | in[55];
assign internal[150] = in[42] ^ in[66];
assign internal[151] = ~(in[49] & in[77] & in[91]);
assign internal[152] = in[56] & in[88];
assign internal[153] = in[63] | in[99];
assign internal[154] = in[70] ^ in[110];
assign internal[155] = ~(in[77] & in[121] & in[143]);
assign internal[156] = in[84] & in[132];
assign internal[157] = in[91] | in[143];
assign internal[158] = in[98] ^ in[10];
assign internal[159] = ~(in[105] & in[21] & in[51]);
assign internal[160] = in[112] & in[32];
assign internal[161] = in[119] | in[43];
assign internal[162] = in[126] ^ in[54];
assign internal[163] = ~(in[133] & in[65] & in[103]);
assign internal[164] = in[140] & in[76];
assign internal[165] = in[3] | in[87];
assign internal[166] = in[10] ^ in[98];
assign internal[167] = ~(in[17] & in[109] & in[11]);
assign internal[168] = in[24] & in[120];
assign internal[169] = in[31] | in[131];
assign internal[170] = in[38] ^ in[142];
assign internal[171] = ~(in[45] & in[9] & in[63]);
assign internal[172] = in[52] & in[20];
assign internal[173] = in[59] | in[31];
assign internal[174] = in[66] ^ in[42];
assign internal[175] = ~(in[73] & in[53] & in[115]);
assign internal[176] = in[80] & in[64];
assign internal[177] = in[87] | in[75];
assign internal[178] = in[94] ^ in[86];
assign internal[179] = ~(in[101] & in[97] & in[23]);
assign internal[180] = in[108] & in[108];
assign internal[181] = in[115] | in[119];
assign internal[182] = in[122] ^ in[130];
assign internal[183] = ~(in[129] & in[141] & in[75]);
assign internal[184] = in[136] & in[8];
assign internal[185] = in[143] | in[19];
assign internal[186] = in[6] ^ in[30];
assign internal[187] = ~(in[13] & in[41] & in[127]);
assign internal[188] = in[20] & in[52];
assign internal[189] = in[27] | in[63];
assign internal[190] = in[34] ^ in[74];
assign internal[191] = ~(in[41] & in[85] & in[35]);
assign internal[192] = in[48] & in[96];
assign internal[193] = in[55] | in[107];
assign internal[194] = in[62] ^ in[118];
assign internal[195] = ~(in[69] & in[129] & in[87]);
assign internal[196] = in[76] & in[140];
assign internal[197] = in[83] | in[7];
assign internal[198] = in[90] ^ in[18];
assign internal[199] = ~(in[97] & in[29] & in[139]);
assign internal[200] = in[104] & in[40];
assign internal[201] = in[111] | in[51];
assign internal[202] = in[118] ^ in[62];
assign internal[203] = ~(in[125] & in[73] & in[47]);
assign internal[204] = in[132] & in[84];
assign internal[205] = in[139] | in[95];
assign internal[206] = in[2] ^ in[106];
assign internal[207] = ~(in[9] & in[117] & in[99]);
assign internal[208] = in[16] & in[128];
assign internal[209] = in[23] | in[139];
assign internal[210] = in[30] ^ in[6];
assign internal[211] = ~(in[37] & in[17] & in[7]);
assign internal[212] = in[44] & in[28];
assign internal[213] = in[51] | in[39];
assign internal[214] = in[58] ^ in[50];
assign internal[215] = ~(in[65] & in[61] & in[59]);
assign internal[216] = in[72] & in[72];
assign internal[217] = in[79] | in[83];
assign internal[218] = in[86] ^ in[94];
assign internal[219] = ~(in[93] & in[105] & in[111]);
assign internal[220] = in[100] & in[116];
assign internal[221] = in[107] | in[127];
assign internal[222] = in[114] ^ in[138];
assign internal[223] = ~(in[121] & in[5] & in[19]);
assign internal[224] = in[128] & in[16];
assign internal[225] = in[135] | in[27];
assign internal[226] = in[142] ^ in[38];
assign internal[227] = ~(in[5] & in[49] & in[71]);
assign internal[228] = in[12] & in[60];
assign internal[229] = in[19] | in[71];
assign internal[230] = in[26] ^ in[82];
assign internal[231] = ~(in[33] & in[93] & in[123]);
assign internal[232] = in[40] & in[104];
assign internal[233] = in[47] | in[115];
assign internal[234] = in[54] ^ in[126];
assign internal[235] = ~(in[61] & in[137] & in[31]);
assign internal[236] = in[68] & in[4];
assign internal[237] = in[75] | in[15];
assign internal[238] = in[82] ^ in[26];
assign internal[239] = ~(in[89] & in[37] & in[83]);
assign internal[240] = in[96] & in[48];
assign internal[241] = in[103] | in[59];
assign internal[242] = in[110] ^ in[70];
assign internal[243] = ~(in[117] & in[81] & in[135]);
assign internal[244] = in[124] & in[92];
assign internal[245] = in[131] | in[103];
assign internal[246] = in[138] ^ in[114];
assign internal[247] = ~(in[1] & in[125] & in[43]);
assign internal[248] = in[8] & in[136];
assign internal[249] = in[15] | in[3];
assign internal[250] = in[22] ^ in[14];
assign internal[251] = ~(in[29] & in[25] & in[95]);
assign internal[252] = in[36] & in[36];
assign internal[253] = in[43] | in[47];
assign internal[254] = in[50] ^ in[58];
assign internal[255] = ~(in[57] & in[69] & in[3]);
assign internal[256] = in[64] & in[80];
assign internal[257] = in[71] | in[91];
assign internal[258] = in[78] ^ in[102];
assign internal[259] = ~(in[85] & in[113] & in[55]);
assign internal[260] = in[92] & in[124];
assign internal[261] = in[99] | in[135];
assign internal[262] = in[106] ^ in[2];
assign internal[263] = ~(in[113] & in[13] & in[107]);
assign internal[264] = in[120] & in[24];
assign internal[265] = in[127] | in[35];
assign internal[266] = in[134] ^ in[46];
assign internal[267] = ~(in[141] & in[57] & in[15]);
assign internal[268] = in[4] & in[68];
assign internal[269] = in[11] | in[79];
assign internal[270] = in[18] ^ in[90];
assign internal[271] = ~(in[25] & in[101] & in[67]);
assign internal[272] = in[32] & in[112];
assign internal[273] = in[39] | in[123];
assign internal[274] = in[46] ^ in[134];
assign internal[275] = ~(in[53] & in[1] & in[119]);
assign internal[276] = in[60] & in[12];
assign internal[277] = in[67] | in[23];
assign internal[278] = in[74] ^ in[34];
assign internal[279] = ~(in[81] & in[45] & in[27]);
assign internal[280] = in[88] & in[56];
assign internal[281] = in[95] | in[67];
assign internal[282] = in[102] ^ in[78];
assign internal[283] = ~(in[109] & in[89] & in[79]);
assign internal[284] = in[116] & in[100];
assign internal[285] = in[123] | in[111];
assign internal[286] = in[130] ^ in[122];
assign internal[287] = ~(in[137] & in[133] & in[131]);

assign out[0] = internal[0] & internal[0];
assign out[1] = internal[3] | internal[5];
assign out[2] = internal[6] ^ internal[10] ^ internal[14];
assign out[3] = internal[9] & internal[15];
assign out[4] = internal[12] | internal[20];
assign out[5] = internal[15] ^ internal[25] ^ internal[35];
assign out[6] = internal[18] & internal[30];
assign out[7] = internal[21] | internal[35];
assign out[8] = internal[24] ^ internal[40] ^ internal[56];
assign out[9] = internal[27] & internal[45];
assign out[10] = internal[30] | internal[50];
assign out[11] = internal[33] ^ internal[55] ^ internal[77];
assign out[12] = internal[36] & internal[60];
assign out[13] = internal[39] | internal[65];
assign out[14] = internal[42] ^ internal[70] ^ internal[98];
assign out[15] = internal[45] & internal[75];
assign out[16] = internal[48] | internal[80];
assign out[17] = internal[51] ^ internal[85] ^ internal[119];
assign out[18] = internal[54] & internal[90];
assign out[19] = internal[57] | internal[95];
assign out[20] = internal[60] ^ internal[100] ^ internal[140];
assign out[21] = internal[63] & internal[105];
assign out[22] = internal[66] | internal[110];
assign out[23] = internal[69] ^ internal[115] ^ internal[161];
assign out[24] = internal[72] & internal[120];
assign out[25] = internal[75] | internal[125];
assign out[26] = internal[78] ^ internal[130] ^ internal[182];
assign out[27] = internal[81] & internal[135];
assign out[28] = internal[84] | internal[140];
assign out[29] = internal[87] ^ internal[145] ^ internal[203];
assign out[30] = internal[90] & internal[150];
assign out[31] = internal[93] | internal[155];
assign out[32] = internal[96] ^ internal[160] ^ internal[224];
assign out[33] = internal[99] & internal[165];
assign out[34] = internal[102] | internal[170];
assign out[35] = internal[105] ^ internal[175] ^ internal[245];
assign out[36] = internal[108] & internal[180];
assign out[37] = internal[111] | internal[185];
assign out[38] = internal[114] ^ internal[190] ^ internal[266];
assign out[39] = internal[117] & internal[195];
assign out[40] = internal[120] | internal[200];
assign out[41] = internal[123] ^ internal[205] ^ internal[287];
assign out[42] = internal[126] & internal[210];
assign out[43] = internal[129] | internal[215];
assign out[44] = internal[132] ^ internal[220] ^ internal[20];
assign out[45] = internal[135] & internal[225];
assign out[46] = internal[138] | internal[230];
assign out[47] = internal[141] ^ internal[235] ^ internal[41];
assign out[48] = internal[144] & internal[240];
assign out[49] = internal[147] | internal[245];
assign out[50] = internal[150] ^ internal[250] ^ internal[62];
assign out[51] = internal[153] & internal[255];
assign out[52] = internal[156] | internal[260];
assign out[53] = internal[159] ^ internal[265] ^ internal[83];
assign out[54] = internal[162] & internal[270];
assign out[55] = internal[165] | internal[275];
assign out[56] = internal[168] ^ internal[280] ^ internal[104];
assign out[57] = internal[171] & internal[285];
assign out[58] = internal[174] | internal[2];
assign out[59] = internal[177] ^ internal[7] ^ internal[125];
assign out[60] = internal[180] & internal[12];
assign out[61] = internal[183] | internal[17];
assign out[62] = internal[186] ^ internal[22] ^ internal[146];
assign out[63] = internal[189] & internal[27];
assign out[64] = internal[192] | internal[32];
assign out[65] = internal[195] ^ internal[37] ^ internal[167];
assign out[66] = internal[198] & internal[42];
assign out[67] = internal[201] | internal[47];
assign out[68] = internal[204] ^ internal[52] ^ internal[188];
assign out[69] = internal[207] & internal[57];
assign out[70] = internal[210] | internal[62];
assign out[71] = internal[213] ^ internal[67] ^ internal[209];

endmodule