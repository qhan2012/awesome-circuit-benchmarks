module aig_mix_8_vl8(
    input [175:0] in,
    output [87:0] out
);

// Mixed AIG logic with various patterns
wire [351:0] internal;

assign internal[0] = in[0] & in[0];
assign internal[1] = in[7] | in[11];
assign internal[2] = in[14] ^ in[22];
assign internal[3] = ~(in[21] & in[33] & in[39]);
assign internal[4] = in[28] & in[44];
assign internal[5] = in[35] | in[55];
assign internal[6] = in[42] ^ in[66];
assign internal[7] = ~(in[49] & in[77] & in[91]);
assign internal[8] = in[56] & in[88];
assign internal[9] = in[63] | in[99];
assign internal[10] = in[70] ^ in[110];
assign internal[11] = ~(in[77] & in[121] & in[143]);
assign internal[12] = in[84] & in[132];
assign internal[13] = in[91] | in[143];
assign internal[14] = in[98] ^ in[154];
assign internal[15] = ~(in[105] & in[165] & in[19]);
assign internal[16] = in[112] & in[0];
assign internal[17] = in[119] | in[11];
assign internal[18] = in[126] ^ in[22];
assign internal[19] = ~(in[133] & in[33] & in[71]);
assign internal[20] = in[140] & in[44];
assign internal[21] = in[147] | in[55];
assign internal[22] = in[154] ^ in[66];
assign internal[23] = ~(in[161] & in[77] & in[123]);
assign internal[24] = in[168] & in[88];
assign internal[25] = in[175] | in[99];
assign internal[26] = in[6] ^ in[110];
assign internal[27] = ~(in[13] & in[121] & in[175]);
assign internal[28] = in[20] & in[132];
assign internal[29] = in[27] | in[143];
assign internal[30] = in[34] ^ in[154];
assign internal[31] = ~(in[41] & in[165] & in[51]);
assign internal[32] = in[48] & in[0];
assign internal[33] = in[55] | in[11];
assign internal[34] = in[62] ^ in[22];
assign internal[35] = ~(in[69] & in[33] & in[103]);
assign internal[36] = in[76] & in[44];
assign internal[37] = in[83] | in[55];
assign internal[38] = in[90] ^ in[66];
assign internal[39] = ~(in[97] & in[77] & in[155]);
assign internal[40] = in[104] & in[88];
assign internal[41] = in[111] | in[99];
assign internal[42] = in[118] ^ in[110];
assign internal[43] = ~(in[125] & in[121] & in[31]);
assign internal[44] = in[132] & in[132];
assign internal[45] = in[139] | in[143];
assign internal[46] = in[146] ^ in[154];
assign internal[47] = ~(in[153] & in[165] & in[83]);
assign internal[48] = in[160] & in[0];
assign internal[49] = in[167] | in[11];
assign internal[50] = in[174] ^ in[22];
assign internal[51] = ~(in[5] & in[33] & in[135]);
assign internal[52] = in[12] & in[44];
assign internal[53] = in[19] | in[55];
assign internal[54] = in[26] ^ in[66];
assign internal[55] = ~(in[33] & in[77] & in[11]);
assign internal[56] = in[40] & in[88];
assign internal[57] = in[47] | in[99];
assign internal[58] = in[54] ^ in[110];
assign internal[59] = ~(in[61] & in[121] & in[63]);
assign internal[60] = in[68] & in[132];
assign internal[61] = in[75] | in[143];
assign internal[62] = in[82] ^ in[154];
assign internal[63] = ~(in[89] & in[165] & in[115]);
assign internal[64] = in[96] & in[0];
assign internal[65] = in[103] | in[11];
assign internal[66] = in[110] ^ in[22];
assign internal[67] = ~(in[117] & in[33] & in[167]);
assign internal[68] = in[124] & in[44];
assign internal[69] = in[131] | in[55];
assign internal[70] = in[138] ^ in[66];
assign internal[71] = ~(in[145] & in[77] & in[43]);
assign internal[72] = in[152] & in[88];
assign internal[73] = in[159] | in[99];
assign internal[74] = in[166] ^ in[110];
assign internal[75] = ~(in[173] & in[121] & in[95]);
assign internal[76] = in[4] & in[132];
assign internal[77] = in[11] | in[143];
assign internal[78] = in[18] ^ in[154];
assign internal[79] = ~(in[25] & in[165] & in[147]);
assign internal[80] = in[32] & in[0];
assign internal[81] = in[39] | in[11];
assign internal[82] = in[46] ^ in[22];
assign internal[83] = ~(in[53] & in[33] & in[23]);
assign internal[84] = in[60] & in[44];
assign internal[85] = in[67] | in[55];
assign internal[86] = in[74] ^ in[66];
assign internal[87] = ~(in[81] & in[77] & in[75]);
assign internal[88] = in[88] & in[88];
assign internal[89] = in[95] | in[99];
assign internal[90] = in[102] ^ in[110];
assign internal[91] = ~(in[109] & in[121] & in[127]);
assign internal[92] = in[116] & in[132];
assign internal[93] = in[123] | in[143];
assign internal[94] = in[130] ^ in[154];
assign internal[95] = ~(in[137] & in[165] & in[3]);
assign internal[96] = in[144] & in[0];
assign internal[97] = in[151] | in[11];
assign internal[98] = in[158] ^ in[22];
assign internal[99] = ~(in[165] & in[33] & in[55]);
assign internal[100] = in[172] & in[44];
assign internal[101] = in[3] | in[55];
assign internal[102] = in[10] ^ in[66];
assign internal[103] = ~(in[17] & in[77] & in[107]);
assign internal[104] = in[24] & in[88];
assign internal[105] = in[31] | in[99];
assign internal[106] = in[38] ^ in[110];
assign internal[107] = ~(in[45] & in[121] & in[159]);
assign internal[108] = in[52] & in[132];
assign internal[109] = in[59] | in[143];
assign internal[110] = in[66] ^ in[154];
assign internal[111] = ~(in[73] & in[165] & in[35]);
assign internal[112] = in[80] & in[0];
assign internal[113] = in[87] | in[11];
assign internal[114] = in[94] ^ in[22];
assign internal[115] = ~(in[101] & in[33] & in[87]);
assign internal[116] = in[108] & in[44];
assign internal[117] = in[115] | in[55];
assign internal[118] = in[122] ^ in[66];
assign internal[119] = ~(in[129] & in[77] & in[139]);
assign internal[120] = in[136] & in[88];
assign internal[121] = in[143] | in[99];
assign internal[122] = in[150] ^ in[110];
assign internal[123] = ~(in[157] & in[121] & in[15]);
assign internal[124] = in[164] & in[132];
assign internal[125] = in[171] | in[143];
assign internal[126] = in[2] ^ in[154];
assign internal[127] = ~(in[9] & in[165] & in[67]);
assign internal[128] = in[16] & in[0];
assign internal[129] = in[23] | in[11];
assign internal[130] = in[30] ^ in[22];
assign internal[131] = ~(in[37] & in[33] & in[119]);
assign internal[132] = in[44] & in[44];
assign internal[133] = in[51] | in[55];
assign internal[134] = in[58] ^ in[66];
assign internal[135] = ~(in[65] & in[77] & in[171]);
assign internal[136] = in[72] & in[88];
assign internal[137] = in[79] | in[99];
assign internal[138] = in[86] ^ in[110];
assign internal[139] = ~(in[93] & in[121] & in[47]);
assign internal[140] = in[100] & in[132];
assign internal[141] = in[107] | in[143];
assign internal[142] = in[114] ^ in[154];
assign internal[143] = ~(in[121] & in[165] & in[99]);
assign internal[144] = in[128] & in[0];
assign internal[145] = in[135] | in[11];
assign internal[146] = in[142] ^ in[22];
assign internal[147] = ~(in[149] & in[33] & in[151]);
assign internal[148] = in[156] & in[44];
assign internal[149] = in[163] | in[55];
assign internal[150] = in[170] ^ in[66];
assign internal[151] = ~(in[1] & in[77] & in[27]);
assign internal[152] = in[8] & in[88];
assign internal[153] = in[15] | in[99];
assign internal[154] = in[22] ^ in[110];
assign internal[155] = ~(in[29] & in[121] & in[79]);
assign internal[156] = in[36] & in[132];
assign internal[157] = in[43] | in[143];
assign internal[158] = in[50] ^ in[154];
assign internal[159] = ~(in[57] & in[165] & in[131]);
assign internal[160] = in[64] & in[0];
assign internal[161] = in[71] | in[11];
assign internal[162] = in[78] ^ in[22];
assign internal[163] = ~(in[85] & in[33] & in[7]);
assign internal[164] = in[92] & in[44];
assign internal[165] = in[99] | in[55];
assign internal[166] = in[106] ^ in[66];
assign internal[167] = ~(in[113] & in[77] & in[59]);
assign internal[168] = in[120] & in[88];
assign internal[169] = in[127] | in[99];
assign internal[170] = in[134] ^ in[110];
assign internal[171] = ~(in[141] & in[121] & in[111]);
assign internal[172] = in[148] & in[132];
assign internal[173] = in[155] | in[143];
assign internal[174] = in[162] ^ in[154];
assign internal[175] = ~(in[169] & in[165] & in[163]);
assign internal[176] = in[0] & in[0];
assign internal[177] = in[7] | in[11];
assign internal[178] = in[14] ^ in[22];
assign internal[179] = ~(in[21] & in[33] & in[39]);
assign internal[180] = in[28] & in[44];
assign internal[181] = in[35] | in[55];
assign internal[182] = in[42] ^ in[66];
assign internal[183] = ~(in[49] & in[77] & in[91]);
assign internal[184] = in[56] & in[88];
assign internal[185] = in[63] | in[99];
assign internal[186] = in[70] ^ in[110];
assign internal[187] = ~(in[77] & in[121] & in[143]);
assign internal[188] = in[84] & in[132];
assign internal[189] = in[91] | in[143];
assign internal[190] = in[98] ^ in[154];
assign internal[191] = ~(in[105] & in[165] & in[19]);
assign internal[192] = in[112] & in[0];
assign internal[193] = in[119] | in[11];
assign internal[194] = in[126] ^ in[22];
assign internal[195] = ~(in[133] & in[33] & in[71]);
assign internal[196] = in[140] & in[44];
assign internal[197] = in[147] | in[55];
assign internal[198] = in[154] ^ in[66];
assign internal[199] = ~(in[161] & in[77] & in[123]);
assign internal[200] = in[168] & in[88];
assign internal[201] = in[175] | in[99];
assign internal[202] = in[6] ^ in[110];
assign internal[203] = ~(in[13] & in[121] & in[175]);
assign internal[204] = in[20] & in[132];
assign internal[205] = in[27] | in[143];
assign internal[206] = in[34] ^ in[154];
assign internal[207] = ~(in[41] & in[165] & in[51]);
assign internal[208] = in[48] & in[0];
assign internal[209] = in[55] | in[11];
assign internal[210] = in[62] ^ in[22];
assign internal[211] = ~(in[69] & in[33] & in[103]);
assign internal[212] = in[76] & in[44];
assign internal[213] = in[83] | in[55];
assign internal[214] = in[90] ^ in[66];
assign internal[215] = ~(in[97] & in[77] & in[155]);
assign internal[216] = in[104] & in[88];
assign internal[217] = in[111] | in[99];
assign internal[218] = in[118] ^ in[110];
assign internal[219] = ~(in[125] & in[121] & in[31]);
assign internal[220] = in[132] & in[132];
assign internal[221] = in[139] | in[143];
assign internal[222] = in[146] ^ in[154];
assign internal[223] = ~(in[153] & in[165] & in[83]);
assign internal[224] = in[160] & in[0];
assign internal[225] = in[167] | in[11];
assign internal[226] = in[174] ^ in[22];
assign internal[227] = ~(in[5] & in[33] & in[135]);
assign internal[228] = in[12] & in[44];
assign internal[229] = in[19] | in[55];
assign internal[230] = in[26] ^ in[66];
assign internal[231] = ~(in[33] & in[77] & in[11]);
assign internal[232] = in[40] & in[88];
assign internal[233] = in[47] | in[99];
assign internal[234] = in[54] ^ in[110];
assign internal[235] = ~(in[61] & in[121] & in[63]);
assign internal[236] = in[68] & in[132];
assign internal[237] = in[75] | in[143];
assign internal[238] = in[82] ^ in[154];
assign internal[239] = ~(in[89] & in[165] & in[115]);
assign internal[240] = in[96] & in[0];
assign internal[241] = in[103] | in[11];
assign internal[242] = in[110] ^ in[22];
assign internal[243] = ~(in[117] & in[33] & in[167]);
assign internal[244] = in[124] & in[44];
assign internal[245] = in[131] | in[55];
assign internal[246] = in[138] ^ in[66];
assign internal[247] = ~(in[145] & in[77] & in[43]);
assign internal[248] = in[152] & in[88];
assign internal[249] = in[159] | in[99];
assign internal[250] = in[166] ^ in[110];
assign internal[251] = ~(in[173] & in[121] & in[95]);
assign internal[252] = in[4] & in[132];
assign internal[253] = in[11] | in[143];
assign internal[254] = in[18] ^ in[154];
assign internal[255] = ~(in[25] & in[165] & in[147]);
assign internal[256] = in[32] & in[0];
assign internal[257] = in[39] | in[11];
assign internal[258] = in[46] ^ in[22];
assign internal[259] = ~(in[53] & in[33] & in[23]);
assign internal[260] = in[60] & in[44];
assign internal[261] = in[67] | in[55];
assign internal[262] = in[74] ^ in[66];
assign internal[263] = ~(in[81] & in[77] & in[75]);
assign internal[264] = in[88] & in[88];
assign internal[265] = in[95] | in[99];
assign internal[266] = in[102] ^ in[110];
assign internal[267] = ~(in[109] & in[121] & in[127]);
assign internal[268] = in[116] & in[132];
assign internal[269] = in[123] | in[143];
assign internal[270] = in[130] ^ in[154];
assign internal[271] = ~(in[137] & in[165] & in[3]);
assign internal[272] = in[144] & in[0];
assign internal[273] = in[151] | in[11];
assign internal[274] = in[158] ^ in[22];
assign internal[275] = ~(in[165] & in[33] & in[55]);
assign internal[276] = in[172] & in[44];
assign internal[277] = in[3] | in[55];
assign internal[278] = in[10] ^ in[66];
assign internal[279] = ~(in[17] & in[77] & in[107]);
assign internal[280] = in[24] & in[88];
assign internal[281] = in[31] | in[99];
assign internal[282] = in[38] ^ in[110];
assign internal[283] = ~(in[45] & in[121] & in[159]);
assign internal[284] = in[52] & in[132];
assign internal[285] = in[59] | in[143];
assign internal[286] = in[66] ^ in[154];
assign internal[287] = ~(in[73] & in[165] & in[35]);
assign internal[288] = in[80] & in[0];
assign internal[289] = in[87] | in[11];
assign internal[290] = in[94] ^ in[22];
assign internal[291] = ~(in[101] & in[33] & in[87]);
assign internal[292] = in[108] & in[44];
assign internal[293] = in[115] | in[55];
assign internal[294] = in[122] ^ in[66];
assign internal[295] = ~(in[129] & in[77] & in[139]);
assign internal[296] = in[136] & in[88];
assign internal[297] = in[143] | in[99];
assign internal[298] = in[150] ^ in[110];
assign internal[299] = ~(in[157] & in[121] & in[15]);
assign internal[300] = in[164] & in[132];
assign internal[301] = in[171] | in[143];
assign internal[302] = in[2] ^ in[154];
assign internal[303] = ~(in[9] & in[165] & in[67]);
assign internal[304] = in[16] & in[0];
assign internal[305] = in[23] | in[11];
assign internal[306] = in[30] ^ in[22];
assign internal[307] = ~(in[37] & in[33] & in[119]);
assign internal[308] = in[44] & in[44];
assign internal[309] = in[51] | in[55];
assign internal[310] = in[58] ^ in[66];
assign internal[311] = ~(in[65] & in[77] & in[171]);
assign internal[312] = in[72] & in[88];
assign internal[313] = in[79] | in[99];
assign internal[314] = in[86] ^ in[110];
assign internal[315] = ~(in[93] & in[121] & in[47]);
assign internal[316] = in[100] & in[132];
assign internal[317] = in[107] | in[143];
assign internal[318] = in[114] ^ in[154];
assign internal[319] = ~(in[121] & in[165] & in[99]);
assign internal[320] = in[128] & in[0];
assign internal[321] = in[135] | in[11];
assign internal[322] = in[142] ^ in[22];
assign internal[323] = ~(in[149] & in[33] & in[151]);
assign internal[324] = in[156] & in[44];
assign internal[325] = in[163] | in[55];
assign internal[326] = in[170] ^ in[66];
assign internal[327] = ~(in[1] & in[77] & in[27]);
assign internal[328] = in[8] & in[88];
assign internal[329] = in[15] | in[99];
assign internal[330] = in[22] ^ in[110];
assign internal[331] = ~(in[29] & in[121] & in[79]);
assign internal[332] = in[36] & in[132];
assign internal[333] = in[43] | in[143];
assign internal[334] = in[50] ^ in[154];
assign internal[335] = ~(in[57] & in[165] & in[131]);
assign internal[336] = in[64] & in[0];
assign internal[337] = in[71] | in[11];
assign internal[338] = in[78] ^ in[22];
assign internal[339] = ~(in[85] & in[33] & in[7]);
assign internal[340] = in[92] & in[44];
assign internal[341] = in[99] | in[55];
assign internal[342] = in[106] ^ in[66];
assign internal[343] = ~(in[113] & in[77] & in[59]);
assign internal[344] = in[120] & in[88];
assign internal[345] = in[127] | in[99];
assign internal[346] = in[134] ^ in[110];
assign internal[347] = ~(in[141] & in[121] & in[111]);
assign internal[348] = in[148] & in[132];
assign internal[349] = in[155] | in[143];
assign internal[350] = in[162] ^ in[154];
assign internal[351] = ~(in[169] & in[165] & in[163]);

assign out[0] = internal[0] & internal[0];
assign out[1] = internal[3] | internal[5];
assign out[2] = internal[6] ^ internal[10] ^ internal[14];
assign out[3] = internal[9] & internal[15];
assign out[4] = internal[12] | internal[20];
assign out[5] = internal[15] ^ internal[25] ^ internal[35];
assign out[6] = internal[18] & internal[30];
assign out[7] = internal[21] | internal[35];
assign out[8] = internal[24] ^ internal[40] ^ internal[56];
assign out[9] = internal[27] & internal[45];
assign out[10] = internal[30] | internal[50];
assign out[11] = internal[33] ^ internal[55] ^ internal[77];
assign out[12] = internal[36] & internal[60];
assign out[13] = internal[39] | internal[65];
assign out[14] = internal[42] ^ internal[70] ^ internal[98];
assign out[15] = internal[45] & internal[75];
assign out[16] = internal[48] | internal[80];
assign out[17] = internal[51] ^ internal[85] ^ internal[119];
assign out[18] = internal[54] & internal[90];
assign out[19] = internal[57] | internal[95];
assign out[20] = internal[60] ^ internal[100] ^ internal[140];
assign out[21] = internal[63] & internal[105];
assign out[22] = internal[66] | internal[110];
assign out[23] = internal[69] ^ internal[115] ^ internal[161];
assign out[24] = internal[72] & internal[120];
assign out[25] = internal[75] | internal[125];
assign out[26] = internal[78] ^ internal[130] ^ internal[182];
assign out[27] = internal[81] & internal[135];
assign out[28] = internal[84] | internal[140];
assign out[29] = internal[87] ^ internal[145] ^ internal[203];
assign out[30] = internal[90] & internal[150];
assign out[31] = internal[93] | internal[155];
assign out[32] = internal[96] ^ internal[160] ^ internal[224];
assign out[33] = internal[99] & internal[165];
assign out[34] = internal[102] | internal[170];
assign out[35] = internal[105] ^ internal[175] ^ internal[245];
assign out[36] = internal[108] & internal[180];
assign out[37] = internal[111] | internal[185];
assign out[38] = internal[114] ^ internal[190] ^ internal[266];
assign out[39] = internal[117] & internal[195];
assign out[40] = internal[120] | internal[200];
assign out[41] = internal[123] ^ internal[205] ^ internal[287];
assign out[42] = internal[126] & internal[210];
assign out[43] = internal[129] | internal[215];
assign out[44] = internal[132] ^ internal[220] ^ internal[308];
assign out[45] = internal[135] & internal[225];
assign out[46] = internal[138] | internal[230];
assign out[47] = internal[141] ^ internal[235] ^ internal[329];
assign out[48] = internal[144] & internal[240];
assign out[49] = internal[147] | internal[245];
assign out[50] = internal[150] ^ internal[250] ^ internal[350];
assign out[51] = internal[153] & internal[255];
assign out[52] = internal[156] | internal[260];
assign out[53] = internal[159] ^ internal[265] ^ internal[19];
assign out[54] = internal[162] & internal[270];
assign out[55] = internal[165] | internal[275];
assign out[56] = internal[168] ^ internal[280] ^ internal[40];
assign out[57] = internal[171] & internal[285];
assign out[58] = internal[174] | internal[290];
assign out[59] = internal[177] ^ internal[295] ^ internal[61];
assign out[60] = internal[180] & internal[300];
assign out[61] = internal[183] | internal[305];
assign out[62] = internal[186] ^ internal[310] ^ internal[82];
assign out[63] = internal[189] & internal[315];
assign out[64] = internal[192] | internal[320];
assign out[65] = internal[195] ^ internal[325] ^ internal[103];
assign out[66] = internal[198] & internal[330];
assign out[67] = internal[201] | internal[335];
assign out[68] = internal[204] ^ internal[340] ^ internal[124];
assign out[69] = internal[207] & internal[345];
assign out[70] = internal[210] | internal[350];
assign out[71] = internal[213] ^ internal[3] ^ internal[145];
assign out[72] = internal[216] & internal[8];
assign out[73] = internal[219] | internal[13];
assign out[74] = internal[222] ^ internal[18] ^ internal[166];
assign out[75] = internal[225] & internal[23];
assign out[76] = internal[228] | internal[28];
assign out[77] = internal[231] ^ internal[33] ^ internal[187];
assign out[78] = internal[234] & internal[38];
assign out[79] = internal[237] | internal[43];
assign out[80] = internal[240] ^ internal[48] ^ internal[208];
assign out[81] = internal[243] & internal[53];
assign out[82] = internal[246] | internal[58];
assign out[83] = internal[249] ^ internal[63] ^ internal[229];
assign out[84] = internal[252] & internal[68];
assign out[85] = internal[255] | internal[73];
assign out[86] = internal[258] ^ internal[78] ^ internal[250];
assign out[87] = internal[261] & internal[83];

endmodule