module conv_5x5_4ch_vl6(
    input [199:0] pixels_in,          // 25 input pixels (packed)
    output [63:0] result_out      // 4 output channels (packed)
);

// Unpack input pixels
wire [7:0] pixel [24:0];
assign pixel[0] = pixels_in[7:0];
assign pixel[1] = pixels_in[15:8];
assign pixel[2] = pixels_in[23:16];
assign pixel[3] = pixels_in[31:24];
assign pixel[4] = pixels_in[39:32];
assign pixel[5] = pixels_in[47:40];
assign pixel[6] = pixels_in[55:48];
assign pixel[7] = pixels_in[63:56];
assign pixel[8] = pixels_in[71:64];
assign pixel[9] = pixels_in[79:72];
assign pixel[10] = pixels_in[87:80];
assign pixel[11] = pixels_in[95:88];
assign pixel[12] = pixels_in[103:96];
assign pixel[13] = pixels_in[111:104];
assign pixel[14] = pixels_in[119:112];
assign pixel[15] = pixels_in[127:120];
assign pixel[16] = pixels_in[135:128];
assign pixel[17] = pixels_in[143:136];
assign pixel[18] = pixels_in[151:144];
assign pixel[19] = pixels_in[159:152];
assign pixel[20] = pixels_in[167:160];
assign pixel[21] = pixels_in[175:168];
assign pixel[22] = pixels_in[183:176];
assign pixel[23] = pixels_in[191:184];
assign pixel[24] = pixels_in[199:192];

// Convolution weights as parameters
// Channel 0 weights
localparam [7:0] WEIGHT_0_0 = 8'd2;
localparam [7:0] WEIGHT_0_1 = 8'd3;
localparam [7:0] WEIGHT_0_2 = 8'd4;
localparam [7:0] WEIGHT_0_3 = 8'd5;
localparam [7:0] WEIGHT_0_4 = 8'd6;
localparam [7:0] WEIGHT_0_5 = 8'd7;
localparam [7:0] WEIGHT_0_6 = 8'd8;
localparam [7:0] WEIGHT_0_7 = 8'd9;
localparam [7:0] WEIGHT_0_8 = 8'd10;
localparam [7:0] WEIGHT_0_9 = 8'd11;
localparam [7:0] WEIGHT_0_10 = 8'd12;
localparam [7:0] WEIGHT_0_11 = 8'd13;
localparam [7:0] WEIGHT_0_12 = 8'd14;
localparam [7:0] WEIGHT_0_13 = 8'd15;
localparam [7:0] WEIGHT_0_14 = 8'd16;
localparam [7:0] WEIGHT_0_15 = 8'd1;
localparam [7:0] WEIGHT_0_16 = 8'd2;
localparam [7:0] WEIGHT_0_17 = 8'd3;
localparam [7:0] WEIGHT_0_18 = 8'd4;
localparam [7:0] WEIGHT_0_19 = 8'd5;
localparam [7:0] WEIGHT_0_20 = 8'd6;
localparam [7:0] WEIGHT_0_21 = 8'd7;
localparam [7:0] WEIGHT_0_22 = 8'd8;
localparam [7:0] WEIGHT_0_23 = 8'd9;
localparam [7:0] WEIGHT_0_24 = 8'd10;
// Channel 1 weights
localparam [7:0] WEIGHT_1_0 = 8'd3;
localparam [7:0] WEIGHT_1_1 = 8'd4;
localparam [7:0] WEIGHT_1_2 = 8'd5;
localparam [7:0] WEIGHT_1_3 = 8'd6;
localparam [7:0] WEIGHT_1_4 = 8'd7;
localparam [7:0] WEIGHT_1_5 = 8'd8;
localparam [7:0] WEIGHT_1_6 = 8'd9;
localparam [7:0] WEIGHT_1_7 = 8'd10;
localparam [7:0] WEIGHT_1_8 = 8'd11;
localparam [7:0] WEIGHT_1_9 = 8'd12;
localparam [7:0] WEIGHT_1_10 = 8'd13;
localparam [7:0] WEIGHT_1_11 = 8'd14;
localparam [7:0] WEIGHT_1_12 = 8'd15;
localparam [7:0] WEIGHT_1_13 = 8'd16;
localparam [7:0] WEIGHT_1_14 = 8'd1;
localparam [7:0] WEIGHT_1_15 = 8'd2;
localparam [7:0] WEIGHT_1_16 = 8'd3;
localparam [7:0] WEIGHT_1_17 = 8'd4;
localparam [7:0] WEIGHT_1_18 = 8'd5;
localparam [7:0] WEIGHT_1_19 = 8'd6;
localparam [7:0] WEIGHT_1_20 = 8'd7;
localparam [7:0] WEIGHT_1_21 = 8'd8;
localparam [7:0] WEIGHT_1_22 = 8'd9;
localparam [7:0] WEIGHT_1_23 = 8'd10;
localparam [7:0] WEIGHT_1_24 = 8'd11;
// Channel 2 weights
localparam [7:0] WEIGHT_2_0 = 8'd4;
localparam [7:0] WEIGHT_2_1 = 8'd5;
localparam [7:0] WEIGHT_2_2 = 8'd6;
localparam [7:0] WEIGHT_2_3 = 8'd7;
localparam [7:0] WEIGHT_2_4 = 8'd8;
localparam [7:0] WEIGHT_2_5 = 8'd9;
localparam [7:0] WEIGHT_2_6 = 8'd10;
localparam [7:0] WEIGHT_2_7 = 8'd11;
localparam [7:0] WEIGHT_2_8 = 8'd12;
localparam [7:0] WEIGHT_2_9 = 8'd13;
localparam [7:0] WEIGHT_2_10 = 8'd14;
localparam [7:0] WEIGHT_2_11 = 8'd15;
localparam [7:0] WEIGHT_2_12 = 8'd16;
localparam [7:0] WEIGHT_2_13 = 8'd1;
localparam [7:0] WEIGHT_2_14 = 8'd2;
localparam [7:0] WEIGHT_2_15 = 8'd3;
localparam [7:0] WEIGHT_2_16 = 8'd4;
localparam [7:0] WEIGHT_2_17 = 8'd5;
localparam [7:0] WEIGHT_2_18 = 8'd6;
localparam [7:0] WEIGHT_2_19 = 8'd7;
localparam [7:0] WEIGHT_2_20 = 8'd8;
localparam [7:0] WEIGHT_2_21 = 8'd9;
localparam [7:0] WEIGHT_2_22 = 8'd10;
localparam [7:0] WEIGHT_2_23 = 8'd11;
localparam [7:0] WEIGHT_2_24 = 8'd12;
// Channel 3 weights
localparam [7:0] WEIGHT_3_0 = 8'd5;
localparam [7:0] WEIGHT_3_1 = 8'd6;
localparam [7:0] WEIGHT_3_2 = 8'd7;
localparam [7:0] WEIGHT_3_3 = 8'd8;
localparam [7:0] WEIGHT_3_4 = 8'd9;
localparam [7:0] WEIGHT_3_5 = 8'd10;
localparam [7:0] WEIGHT_3_6 = 8'd11;
localparam [7:0] WEIGHT_3_7 = 8'd12;
localparam [7:0] WEIGHT_3_8 = 8'd13;
localparam [7:0] WEIGHT_3_9 = 8'd14;
localparam [7:0] WEIGHT_3_10 = 8'd15;
localparam [7:0] WEIGHT_3_11 = 8'd16;
localparam [7:0] WEIGHT_3_12 = 8'd1;
localparam [7:0] WEIGHT_3_13 = 8'd2;
localparam [7:0] WEIGHT_3_14 = 8'd3;
localparam [7:0] WEIGHT_3_15 = 8'd4;
localparam [7:0] WEIGHT_3_16 = 8'd5;
localparam [7:0] WEIGHT_3_17 = 8'd6;
localparam [7:0] WEIGHT_3_18 = 8'd7;
localparam [7:0] WEIGHT_3_19 = 8'd8;
localparam [7:0] WEIGHT_3_20 = 8'd9;
localparam [7:0] WEIGHT_3_21 = 8'd10;
localparam [7:0] WEIGHT_3_22 = 8'd11;
localparam [7:0] WEIGHT_3_23 = 8'd12;
localparam [7:0] WEIGHT_3_24 = 8'd13;

// Output channels
wire [15:0] channel_out [3:0];

// Parallel convolution computation for each channel
// Channel 0 computation
wire [15:0] products_0 [24:0];
assign products_0[0] = pixel[0] * WEIGHT_0_0;
assign products_0[1] = pixel[1] * WEIGHT_0_1;
assign products_0[2] = pixel[2] * WEIGHT_0_2;
assign products_0[3] = pixel[3] * WEIGHT_0_3;
assign products_0[4] = pixel[4] * WEIGHT_0_4;
assign products_0[5] = pixel[5] * WEIGHT_0_5;
assign products_0[6] = pixel[6] * WEIGHT_0_6;
assign products_0[7] = pixel[7] * WEIGHT_0_7;
assign products_0[8] = pixel[8] * WEIGHT_0_8;
assign products_0[9] = pixel[9] * WEIGHT_0_9;
assign products_0[10] = pixel[10] * WEIGHT_0_10;
assign products_0[11] = pixel[11] * WEIGHT_0_11;
assign products_0[12] = pixel[12] * WEIGHT_0_12;
assign products_0[13] = pixel[13] * WEIGHT_0_13;
assign products_0[14] = pixel[14] * WEIGHT_0_14;
assign products_0[15] = pixel[15] * WEIGHT_0_15;
assign products_0[16] = pixel[16] * WEIGHT_0_16;
assign products_0[17] = pixel[17] * WEIGHT_0_17;
assign products_0[18] = pixel[18] * WEIGHT_0_18;
assign products_0[19] = pixel[19] * WEIGHT_0_19;
assign products_0[20] = pixel[20] * WEIGHT_0_20;
assign products_0[21] = pixel[21] * WEIGHT_0_21;
assign products_0[22] = pixel[22] * WEIGHT_0_22;
assign products_0[23] = pixel[23] * WEIGHT_0_23;
assign products_0[24] = pixel[24] * WEIGHT_0_24;
assign channel_out[0] = products_0[0] + products_0[1] + products_0[2] + products_0[3] + products_0[4] + products_0[5] + products_0[6] + products_0[7] + products_0[8] + products_0[9] + products_0[10] + products_0[11] + products_0[12] + products_0[13] + products_0[14] + products_0[15] + products_0[16] + products_0[17] + products_0[18] + products_0[19] + products_0[20] + products_0[21] + products_0[22] + products_0[23] + products_0[24];
// Channel 1 computation
wire [15:0] products_1 [24:0];
assign products_1[0] = pixel[0] * WEIGHT_1_0;
assign products_1[1] = pixel[1] * WEIGHT_1_1;
assign products_1[2] = pixel[2] * WEIGHT_1_2;
assign products_1[3] = pixel[3] * WEIGHT_1_3;
assign products_1[4] = pixel[4] * WEIGHT_1_4;
assign products_1[5] = pixel[5] * WEIGHT_1_5;
assign products_1[6] = pixel[6] * WEIGHT_1_6;
assign products_1[7] = pixel[7] * WEIGHT_1_7;
assign products_1[8] = pixel[8] * WEIGHT_1_8;
assign products_1[9] = pixel[9] * WEIGHT_1_9;
assign products_1[10] = pixel[10] * WEIGHT_1_10;
assign products_1[11] = pixel[11] * WEIGHT_1_11;
assign products_1[12] = pixel[12] * WEIGHT_1_12;
assign products_1[13] = pixel[13] * WEIGHT_1_13;
assign products_1[14] = pixel[14] * WEIGHT_1_14;
assign products_1[15] = pixel[15] * WEIGHT_1_15;
assign products_1[16] = pixel[16] * WEIGHT_1_16;
assign products_1[17] = pixel[17] * WEIGHT_1_17;
assign products_1[18] = pixel[18] * WEIGHT_1_18;
assign products_1[19] = pixel[19] * WEIGHT_1_19;
assign products_1[20] = pixel[20] * WEIGHT_1_20;
assign products_1[21] = pixel[21] * WEIGHT_1_21;
assign products_1[22] = pixel[22] * WEIGHT_1_22;
assign products_1[23] = pixel[23] * WEIGHT_1_23;
assign products_1[24] = pixel[24] * WEIGHT_1_24;
assign channel_out[1] = products_1[0] + products_1[1] + products_1[2] + products_1[3] + products_1[4] + products_1[5] + products_1[6] + products_1[7] + products_1[8] + products_1[9] + products_1[10] + products_1[11] + products_1[12] + products_1[13] + products_1[14] + products_1[15] + products_1[16] + products_1[17] + products_1[18] + products_1[19] + products_1[20] + products_1[21] + products_1[22] + products_1[23] + products_1[24];
// Channel 2 computation
wire [15:0] products_2 [24:0];
assign products_2[0] = pixel[0] * WEIGHT_2_0;
assign products_2[1] = pixel[1] * WEIGHT_2_1;
assign products_2[2] = pixel[2] * WEIGHT_2_2;
assign products_2[3] = pixel[3] * WEIGHT_2_3;
assign products_2[4] = pixel[4] * WEIGHT_2_4;
assign products_2[5] = pixel[5] * WEIGHT_2_5;
assign products_2[6] = pixel[6] * WEIGHT_2_6;
assign products_2[7] = pixel[7] * WEIGHT_2_7;
assign products_2[8] = pixel[8] * WEIGHT_2_8;
assign products_2[9] = pixel[9] * WEIGHT_2_9;
assign products_2[10] = pixel[10] * WEIGHT_2_10;
assign products_2[11] = pixel[11] * WEIGHT_2_11;
assign products_2[12] = pixel[12] * WEIGHT_2_12;
assign products_2[13] = pixel[13] * WEIGHT_2_13;
assign products_2[14] = pixel[14] * WEIGHT_2_14;
assign products_2[15] = pixel[15] * WEIGHT_2_15;
assign products_2[16] = pixel[16] * WEIGHT_2_16;
assign products_2[17] = pixel[17] * WEIGHT_2_17;
assign products_2[18] = pixel[18] * WEIGHT_2_18;
assign products_2[19] = pixel[19] * WEIGHT_2_19;
assign products_2[20] = pixel[20] * WEIGHT_2_20;
assign products_2[21] = pixel[21] * WEIGHT_2_21;
assign products_2[22] = pixel[22] * WEIGHT_2_22;
assign products_2[23] = pixel[23] * WEIGHT_2_23;
assign products_2[24] = pixel[24] * WEIGHT_2_24;
assign channel_out[2] = products_2[0] + products_2[1] + products_2[2] + products_2[3] + products_2[4] + products_2[5] + products_2[6] + products_2[7] + products_2[8] + products_2[9] + products_2[10] + products_2[11] + products_2[12] + products_2[13] + products_2[14] + products_2[15] + products_2[16] + products_2[17] + products_2[18] + products_2[19] + products_2[20] + products_2[21] + products_2[22] + products_2[23] + products_2[24];
// Channel 3 computation
wire [15:0] products_3 [24:0];
assign products_3[0] = pixel[0] * WEIGHT_3_0;
assign products_3[1] = pixel[1] * WEIGHT_3_1;
assign products_3[2] = pixel[2] * WEIGHT_3_2;
assign products_3[3] = pixel[3] * WEIGHT_3_3;
assign products_3[4] = pixel[4] * WEIGHT_3_4;
assign products_3[5] = pixel[5] * WEIGHT_3_5;
assign products_3[6] = pixel[6] * WEIGHT_3_6;
assign products_3[7] = pixel[7] * WEIGHT_3_7;
assign products_3[8] = pixel[8] * WEIGHT_3_8;
assign products_3[9] = pixel[9] * WEIGHT_3_9;
assign products_3[10] = pixel[10] * WEIGHT_3_10;
assign products_3[11] = pixel[11] * WEIGHT_3_11;
assign products_3[12] = pixel[12] * WEIGHT_3_12;
assign products_3[13] = pixel[13] * WEIGHT_3_13;
assign products_3[14] = pixel[14] * WEIGHT_3_14;
assign products_3[15] = pixel[15] * WEIGHT_3_15;
assign products_3[16] = pixel[16] * WEIGHT_3_16;
assign products_3[17] = pixel[17] * WEIGHT_3_17;
assign products_3[18] = pixel[18] * WEIGHT_3_18;
assign products_3[19] = pixel[19] * WEIGHT_3_19;
assign products_3[20] = pixel[20] * WEIGHT_3_20;
assign products_3[21] = pixel[21] * WEIGHT_3_21;
assign products_3[22] = pixel[22] * WEIGHT_3_22;
assign products_3[23] = pixel[23] * WEIGHT_3_23;
assign products_3[24] = pixel[24] * WEIGHT_3_24;
assign channel_out[3] = products_3[0] + products_3[1] + products_3[2] + products_3[3] + products_3[4] + products_3[5] + products_3[6] + products_3[7] + products_3[8] + products_3[9] + products_3[10] + products_3[11] + products_3[12] + products_3[13] + products_3[14] + products_3[15] + products_3[16] + products_3[17] + products_3[18] + products_3[19] + products_3[20] + products_3[21] + products_3[22] + products_3[23] + products_3[24];

// Pack output channels
assign result_out[15:0] = channel_out[0];
assign result_out[31:16] = channel_out[1];
assign result_out[47:32] = channel_out[2];
assign result_out[63:48] = channel_out[3];

endmodule