module mult_8x8_dadda_l4(
    input [7:0] a,
    input [7:0] b,
    output [15:0] product
);

// Wallace tree multiplier (simplified)
wire [63:0] pp;

// Generate partial products
genvar i, j;
generate
    for (i = 0; i < 8; i = i + 1) begin: pp_row
        for (j = 0; j < 8; j = j + 1) begin: pp_col
            assign pp[i*8+j] = a[j] & b[i];
        end
    end
endgenerate

// Wallace tree reduction (simplified - actual implementation would be more complex)
reg [15:0] sum;
integer k, l;
always @(*) begin
    sum = 16'b0;
    for (k = 0; k < 8; k = k + 1) begin
        for (l = 0; l < 8; l = l + 1) begin
            sum = sum + (pp[k*8+l] << (k+l));
        end
    end
end

assign product = sum;

endmodule