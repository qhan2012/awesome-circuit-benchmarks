module aig_mix_2_vl2(
    input [79:0] in,
    output [39:0] out
);

// Mixed AIG logic with various patterns
wire [159:0] internal;

assign internal[0] = in[0] & in[0];
assign internal[1] = in[7] | in[11];
assign internal[2] = in[14] ^ in[22];
assign internal[3] = ~(in[21] & in[33] & in[39]);
assign internal[4] = in[28] & in[44];
assign internal[5] = in[35] | in[55];
assign internal[6] = in[42] ^ in[66];
assign internal[7] = ~(in[49] & in[77] & in[11]);
assign internal[8] = in[56] & in[8];
assign internal[9] = in[63] | in[19];
assign internal[10] = in[70] ^ in[30];
assign internal[11] = ~(in[77] & in[41] & in[63]);
assign internal[12] = in[4] & in[52];
assign internal[13] = in[11] | in[63];
assign internal[14] = in[18] ^ in[74];
assign internal[15] = ~(in[25] & in[5] & in[35]);
assign internal[16] = in[32] & in[16];
assign internal[17] = in[39] | in[27];
assign internal[18] = in[46] ^ in[38];
assign internal[19] = ~(in[53] & in[49] & in[7]);
assign internal[20] = in[60] & in[60];
assign internal[21] = in[67] | in[71];
assign internal[22] = in[74] ^ in[2];
assign internal[23] = ~(in[1] & in[13] & in[59]);
assign internal[24] = in[8] & in[24];
assign internal[25] = in[15] | in[35];
assign internal[26] = in[22] ^ in[46];
assign internal[27] = ~(in[29] & in[57] & in[31]);
assign internal[28] = in[36] & in[68];
assign internal[29] = in[43] | in[79];
assign internal[30] = in[50] ^ in[10];
assign internal[31] = ~(in[57] & in[21] & in[3]);
assign internal[32] = in[64] & in[32];
assign internal[33] = in[71] | in[43];
assign internal[34] = in[78] ^ in[54];
assign internal[35] = ~(in[5] & in[65] & in[55]);
assign internal[36] = in[12] & in[76];
assign internal[37] = in[19] | in[7];
assign internal[38] = in[26] ^ in[18];
assign internal[39] = ~(in[33] & in[29] & in[27]);
assign internal[40] = in[40] & in[40];
assign internal[41] = in[47] | in[51];
assign internal[42] = in[54] ^ in[62];
assign internal[43] = ~(in[61] & in[73] & in[79]);
assign internal[44] = in[68] & in[4];
assign internal[45] = in[75] | in[15];
assign internal[46] = in[2] ^ in[26];
assign internal[47] = ~(in[9] & in[37] & in[51]);
assign internal[48] = in[16] & in[48];
assign internal[49] = in[23] | in[59];
assign internal[50] = in[30] ^ in[70];
assign internal[51] = ~(in[37] & in[1] & in[23]);
assign internal[52] = in[44] & in[12];
assign internal[53] = in[51] | in[23];
assign internal[54] = in[58] ^ in[34];
assign internal[55] = ~(in[65] & in[45] & in[75]);
assign internal[56] = in[72] & in[56];
assign internal[57] = in[79] | in[67];
assign internal[58] = in[6] ^ in[78];
assign internal[59] = ~(in[13] & in[9] & in[47]);
assign internal[60] = in[20] & in[20];
assign internal[61] = in[27] | in[31];
assign internal[62] = in[34] ^ in[42];
assign internal[63] = ~(in[41] & in[53] & in[19]);
assign internal[64] = in[48] & in[64];
assign internal[65] = in[55] | in[75];
assign internal[66] = in[62] ^ in[6];
assign internal[67] = ~(in[69] & in[17] & in[71]);
assign internal[68] = in[76] & in[28];
assign internal[69] = in[3] | in[39];
assign internal[70] = in[10] ^ in[50];
assign internal[71] = ~(in[17] & in[61] & in[43]);
assign internal[72] = in[24] & in[72];
assign internal[73] = in[31] | in[3];
assign internal[74] = in[38] ^ in[14];
assign internal[75] = ~(in[45] & in[25] & in[15]);
assign internal[76] = in[52] & in[36];
assign internal[77] = in[59] | in[47];
assign internal[78] = in[66] ^ in[58];
assign internal[79] = ~(in[73] & in[69] & in[67]);
assign internal[80] = in[0] & in[0];
assign internal[81] = in[7] | in[11];
assign internal[82] = in[14] ^ in[22];
assign internal[83] = ~(in[21] & in[33] & in[39]);
assign internal[84] = in[28] & in[44];
assign internal[85] = in[35] | in[55];
assign internal[86] = in[42] ^ in[66];
assign internal[87] = ~(in[49] & in[77] & in[11]);
assign internal[88] = in[56] & in[8];
assign internal[89] = in[63] | in[19];
assign internal[90] = in[70] ^ in[30];
assign internal[91] = ~(in[77] & in[41] & in[63]);
assign internal[92] = in[4] & in[52];
assign internal[93] = in[11] | in[63];
assign internal[94] = in[18] ^ in[74];
assign internal[95] = ~(in[25] & in[5] & in[35]);
assign internal[96] = in[32] & in[16];
assign internal[97] = in[39] | in[27];
assign internal[98] = in[46] ^ in[38];
assign internal[99] = ~(in[53] & in[49] & in[7]);
assign internal[100] = in[60] & in[60];
assign internal[101] = in[67] | in[71];
assign internal[102] = in[74] ^ in[2];
assign internal[103] = ~(in[1] & in[13] & in[59]);
assign internal[104] = in[8] & in[24];
assign internal[105] = in[15] | in[35];
assign internal[106] = in[22] ^ in[46];
assign internal[107] = ~(in[29] & in[57] & in[31]);
assign internal[108] = in[36] & in[68];
assign internal[109] = in[43] | in[79];
assign internal[110] = in[50] ^ in[10];
assign internal[111] = ~(in[57] & in[21] & in[3]);
assign internal[112] = in[64] & in[32];
assign internal[113] = in[71] | in[43];
assign internal[114] = in[78] ^ in[54];
assign internal[115] = ~(in[5] & in[65] & in[55]);
assign internal[116] = in[12] & in[76];
assign internal[117] = in[19] | in[7];
assign internal[118] = in[26] ^ in[18];
assign internal[119] = ~(in[33] & in[29] & in[27]);
assign internal[120] = in[40] & in[40];
assign internal[121] = in[47] | in[51];
assign internal[122] = in[54] ^ in[62];
assign internal[123] = ~(in[61] & in[73] & in[79]);
assign internal[124] = in[68] & in[4];
assign internal[125] = in[75] | in[15];
assign internal[126] = in[2] ^ in[26];
assign internal[127] = ~(in[9] & in[37] & in[51]);
assign internal[128] = in[16] & in[48];
assign internal[129] = in[23] | in[59];
assign internal[130] = in[30] ^ in[70];
assign internal[131] = ~(in[37] & in[1] & in[23]);
assign internal[132] = in[44] & in[12];
assign internal[133] = in[51] | in[23];
assign internal[134] = in[58] ^ in[34];
assign internal[135] = ~(in[65] & in[45] & in[75]);
assign internal[136] = in[72] & in[56];
assign internal[137] = in[79] | in[67];
assign internal[138] = in[6] ^ in[78];
assign internal[139] = ~(in[13] & in[9] & in[47]);
assign internal[140] = in[20] & in[20];
assign internal[141] = in[27] | in[31];
assign internal[142] = in[34] ^ in[42];
assign internal[143] = ~(in[41] & in[53] & in[19]);
assign internal[144] = in[48] & in[64];
assign internal[145] = in[55] | in[75];
assign internal[146] = in[62] ^ in[6];
assign internal[147] = ~(in[69] & in[17] & in[71]);
assign internal[148] = in[76] & in[28];
assign internal[149] = in[3] | in[39];
assign internal[150] = in[10] ^ in[50];
assign internal[151] = ~(in[17] & in[61] & in[43]);
assign internal[152] = in[24] & in[72];
assign internal[153] = in[31] | in[3];
assign internal[154] = in[38] ^ in[14];
assign internal[155] = ~(in[45] & in[25] & in[15]);
assign internal[156] = in[52] & in[36];
assign internal[157] = in[59] | in[47];
assign internal[158] = in[66] ^ in[58];
assign internal[159] = ~(in[73] & in[69] & in[67]);

assign out[0] = internal[0] & internal[0];
assign out[1] = internal[3] | internal[5];
assign out[2] = internal[6] ^ internal[10] ^ internal[14];
assign out[3] = internal[9] & internal[15];
assign out[4] = internal[12] | internal[20];
assign out[5] = internal[15] ^ internal[25] ^ internal[35];
assign out[6] = internal[18] & internal[30];
assign out[7] = internal[21] | internal[35];
assign out[8] = internal[24] ^ internal[40] ^ internal[56];
assign out[9] = internal[27] & internal[45];
assign out[10] = internal[30] | internal[50];
assign out[11] = internal[33] ^ internal[55] ^ internal[77];
assign out[12] = internal[36] & internal[60];
assign out[13] = internal[39] | internal[65];
assign out[14] = internal[42] ^ internal[70] ^ internal[98];
assign out[15] = internal[45] & internal[75];
assign out[16] = internal[48] | internal[80];
assign out[17] = internal[51] ^ internal[85] ^ internal[119];
assign out[18] = internal[54] & internal[90];
assign out[19] = internal[57] | internal[95];
assign out[20] = internal[60] ^ internal[100] ^ internal[140];
assign out[21] = internal[63] & internal[105];
assign out[22] = internal[66] | internal[110];
assign out[23] = internal[69] ^ internal[115] ^ internal[1];
assign out[24] = internal[72] & internal[120];
assign out[25] = internal[75] | internal[125];
assign out[26] = internal[78] ^ internal[130] ^ internal[22];
assign out[27] = internal[81] & internal[135];
assign out[28] = internal[84] | internal[140];
assign out[29] = internal[87] ^ internal[145] ^ internal[43];
assign out[30] = internal[90] & internal[150];
assign out[31] = internal[93] | internal[155];
assign out[32] = internal[96] ^ internal[0] ^ internal[64];
assign out[33] = internal[99] & internal[5];
assign out[34] = internal[102] | internal[10];
assign out[35] = internal[105] ^ internal[15] ^ internal[85];
assign out[36] = internal[108] & internal[20];
assign out[37] = internal[111] | internal[25];
assign out[38] = internal[114] ^ internal[30] ^ internal[106];
assign out[39] = internal[117] & internal[35];

endmodule